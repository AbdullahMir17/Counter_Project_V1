//dusfds